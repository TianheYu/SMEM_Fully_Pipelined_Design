`define PER_H 2.5

module sim_RAM_read();
	parameter DONE = 6'b11111;
	
	reg reset_n;
	reg clk;
	reg [5:0] status_read;
	reg [5:0] status_query;
	
	// part 1: load all reads
	reg load_valid;
	reg [511:0] 		load_data;
	wire [8:0] curr_num;
	
	// part 2: provide new read to pipeline
	reg new_read; //indicate RAM to update new_read
	wire new_read_valid;
	wire [8:0] new_read_num; //equal to read_num
	wire [63:0] new_ik_x0, new_ik_x1, new_ik_x2, new_ik_info;
	wire [6:0] new_forward_i;
	
	//part 3: provide new query to queue

	reg [6:0] query_position;
	reg [8:0] query_read_num;
	wire [7:0] new_read_query;
	
	wire [63:0] primary;
	wire [63:0] L2_0, L2_1, L2_2, L2_3;

	RAM_read uut(
		.reset_n(reset_n),
		.clk(clk),
		
		
		// part 1: load all reads
		.status_read(status_read),
		.load_valid(load_valid),
		.load_data(load_data),
		.curr_num(curr_num),
		
		// part 2: provide new read to pipeline
		.status_query(status_query),
		.new_read(new_read), //indicate RAM to update new_read
		.new_read_valid(new_read_valid),
		.new_read_num(new_read_num), //equal to read_num
		.new_ik_x0(new_ik_x0), 
		.new_ik_x1(new_ik_x1), 
		.new_ik_x2(new_ik_x2), 
		.new_ik_info(new_ik_info),
		.new_forward_i(new_forward_i),
		
		//part 3: provide new query to queue
		.query_position(query_position),
		.query_read_num(query_read_num),
		.new_read_query(new_read_query),
		
		//part 4: parameters
		.primary(primary),
		.L2_0(L2_0),
		.L2_1(L2_1),
		.L2_2(L2_2),
		.L2_3(L2_3)
	);
	
	initial forever #`PER_H clk = !clk;
	
	initial begin
	
		reset_n = 0;
		clk = 1;
		status_read = DONE;
		status_query = DONE;
		
		load_valid = 0;
		load_data = 0;
	
		new_read = 0; 
	
		query_position = 0;
		query_read_num = 0;
		
		#`PER_H;#`PER_H;
		#0.1
		#`PER_H;#`PER_H;
		#`PER_H;#`PER_H;
		
		reset_n = 1;
		
		#`PER_H;#`PER_H;
		#`PER_H;#`PER_H;
		
		//test part 1
		
		load_valid = 1;
		
		load_data = 512'h00000203030303020000020002000300010303030301030303030100000200030200020200000003010000010301010302030203020300020302010301000303;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001020203030300030002020302000001020301030000020203020303030303010301020100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		
		load_data = 512'h03020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010103030003030202020003030202020003030202020003030202020003030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		
		load_data = 512'h00000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000300;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001000003000101000003010101000103010101000003020101000003010101000003020101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		
		load_data = 512'h03020203000000020202000302020202000300020202000303020202000303020202000000020202000302020202020303020202000300020202000303020300;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010202020003030202020000030002020003000202000003030202020003010202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		
		load_data = 512'h02020103000202020003030202020003010202020003030202020003010202020103010202020003030202020003030202020003030202020003030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020200030302020200030102020200030302020200030302020200030102020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h01000301010100000301000000000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000300;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000002000102000003010101000003010101000003010101000002010101000003010301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02020200020302020200010302020200010302020200020302020200020302020200020302020200010302020200020302020200020302020200010302020200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003020202000103020202000103020202000103020202000103020202000103020202000103;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02030202000102000102010000020200010002020202000100010101010101000001010201000303010201020102030102020200020300010200020101020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010202030202000100010200020001000102010202030200000101020301020202020203;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h01000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02000303020202000303020202000303020202000303020202000303020202000203020202000202020202000201020202000203020202000203020202000203;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020003030202020003030202020003030202020003030202020003030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h00020200030302020201030202020200000102020200030303020201030302020200030302020303030302000200010302020200000303010200030002020200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003000202000002020201020303020301020303020202000201020200000303000202010302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h00010200030101020001020003010001030101030000000101000000030101010003030101010000030101010000030101010000000101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010200010301030100030101010300000001010103010300010100010301030001030301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h00020000020102020303020102020301020200010102000103010101000301010001030203020200000001010302010101020102020301030003010101010200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010103000101000102010200020003000302030203010102030001030101010003010001;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h02020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003020202000303020202000303020202000303020202000303020202000303020202000303;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010301030002010103;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010100000301010100000301010100000301010100000301010100000301010100000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h03010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h01020202020102020102000100010102000202010100010101000102000001010101020202010100010102010202000202020101020302020101020201020302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003000301000102020200010201010101030002020302020200020302010201030000010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h00030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000301010100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h02020200030302020201030302020200030302020201030302020201030302020201030302020201030302020201030302020201030302020201030302020201;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020200030302020200030302020200030302020200030302020200030302020200000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h02000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020003030202020003030202020003030202020003030202020003030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h03010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000002020201;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h02000303020202000303020202000303020202000003020202000003030202000303020202000303020202000303020202000303020202000303020202000303;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020200030302020200030302020200030302020200030302020200030302020203030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h01010000030101010000030101010000030101010000020101010000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010100000001010100000301010100000301010100000301010100000300010100000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h02030303020300030303000202000003000202000302020200000303020202010302020202020300020002000303020202030300020000000303020203000303;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000020303020002020003030103020003030102020303000001020103030100020003000202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h01030200030101020000030101010300030103010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030102030002000102020202010300000301000100010301030100000301020303010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h03030202020000030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003030202020003030202020003030202020003030202020003030202020003030202020000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h01010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010100000301010101000301010100000301010100000301010100000301010100000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h03030202020003030202020003030202020003030202020003030202020003030202020003000202020003000202020003010202020003030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003030100010101020002000302020302010200030302020200030302020200030302020200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h01010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010101030201020001000300010200000201010100000301010100000301010100000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h02020003030202020003030302020003030202020003030202020200030202020203030202020000030202020003030302020003030202020200030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003020200030302020202030302020202030302020200030302020202030302020202030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h01010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010101000003010101030003000101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01010103010100010103010102010102030101010301020203020203000101000100030302020203010000010201010200030302030100030203020303030002;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010102030101010301030200010301010001010103010103000201020001010301020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h01010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h03020001020301010002020002000201010301030302010002010200000101020200020200020102000101010102000201020201010102020200020100010103;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002010103020301020300010101000203020002010302030002010201020000020200010102;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h03030202020003020202020003020202020003020202020003020202020003020202000303020202000303020202000303020202000303020202000303020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000030302020200030202020200030202020200030302020200030202020200030202020200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h03010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h01010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h03020202000302020202000302020202000302020202030302020200030302020200030302020200030302020200030302020203030202020003030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003020202020003020202020003020202020003020202020003030202020003030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02020003030202020003030202020003030202020003030202020003030202020003030202020003030202020003030202020003030202020003030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003020202000303020202000303020202000303020202000303020202030302020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h01010100000301010100000301010100000301010100000301010100000301040100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h00020302020200020302020200030302020200020302020200020202020200030302020200030302020200020302020200030302020200030302020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002000203020202000203020202000303020202000303020202000203020202000303020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h03010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003000101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h00030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030002000202000303020202000303020202000303020202000303020202000303020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h00030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030002000100000301010101000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h00030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030002000100000301010100000301010100000301010100000301010100000301010100;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h00030302020200030302020200030302020200020302020200030302020200030302020200030302020200030302020200030302020200030302020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030002000202000302020202000303020202000303020202000303020202000303020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h02000303020202000003030202000003020202000303020202000303020202000303020202000303020202000303020202000303020202000303020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020003030202020003030202020003030202020003030202020003030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h01000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02000303020202000003020202000003020202000303020202000303020202000303020202000303020202000303020202000303020202000303020200030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020003020202020003030202020003030202020003020202020003030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h03010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h01010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000030101010000;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010100000301010100000301010100000301010100000301010100000301010100000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe0000000105c961890000000000000001;#`PER_H;#`PER_H;
		load_data = 512'h02000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202000303020202030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020003000202020003030202020003030202020003000202020003010202020003020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h00030302020202030302020200030202020000030202020003030202020200030302020200000302020202030302020202000303020202000303020202000303;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002000303020202000303020202000303020202000303020202000303020202000303020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h00000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010000010101000003010101000003010101000003010101000003010101000003010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h00000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301010100000301;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030002000101000003010101000003010101000003010101000003010101000003010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c500000000b8e1c8c4000000006bfa2fff;#`PER_H;#`PER_H;
		load_data = 512'h03030202020003030202020003030202020003030202020003000202020003020202020003030202020003000202020003030202020003030202020003030202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001030002000200030002020200030202020200030202020200030302020200030302020200;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;
		load_data = 512'h01000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001010000030101010000030101010000030101010000030101010000030101010000030101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02020200030302020200030302020200030202020200030202020203030202020203030202020003030202020003030202020003030202020003030202020003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000003020202000302020202000302020202000302020202000303020202000303020202000302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h01000301010101000301010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003010101000003;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000001000000010101000000010101000001010101000003010101000003010101000003010101;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000006bfa2ffe00000000000000010000000105c96189;#`PER_H;#`PER_H;
		load_data = 512'h02020003030202020003020202020003030202020303020202000303020202000301020202020003030002020003030202020003030202020200030302020202;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000002020200030302020200030302020200030202020200030302010200030302020203030302;#`PER_H;#`PER_H;
		load_data = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d383ea000000000000000010000000000000000;#`PER_H;#`PER_H;
		load_data = 512'h0000000105c9618800000000b8e1c8c3000000006bfa2ffe00000000000000000000000000000001000000004ce798c5000000006bfa2fff00000000b8e1c8c4;#`PER_H;#`PER_H;

		load_valid = 0;
		
		//--------------------------------------
		
		//test part 2
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		
		status_read = 0;
		new_read = 1;
		
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;

		new_read = 0;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		
		new_read = 1;
		#300 //60 cycles
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		
		new_read = 0;
		
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		
		// test part 3
		status_read = DONE;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		
		status_query = 0;
		query_read_num = 0; query_position = 0;#`PER_H;	#`PER_H;
		query_read_num = 0; query_position = 1;#`PER_H;	#`PER_H;
		query_read_num = 0; query_position = 2;#`PER_H;	#`PER_H;
		query_read_num = 0; query_position = 3;#`PER_H;	#`PER_H;
		query_read_num = 1; query_position = 0;#`PER_H;	#`PER_H;
		query_read_num = 1; query_position = 1;#`PER_H;	#`PER_H;
		query_read_num = 1; query_position = 2;#`PER_H;	#`PER_H;
		query_read_num = 1; query_position = 3;#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		#`PER_H;	#`PER_H;
		status_query = DONE;
		#`PER_H;	#`PER_H;
		
		
		
		
		$finish;
		
	end
endmodule